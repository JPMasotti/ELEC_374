`timescale 1ns/10ps

module ldi_tb;

endmodule