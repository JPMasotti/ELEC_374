module inport(
    input wire clk, clear,
    input wire [31:0] d,
    output reg [31:0] q
);

  always @(posedge clk) begin
    if (clear)
      q <= 32'b0;
    else
      q <= d;      
  end

endmodule
