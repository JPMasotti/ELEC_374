`timescale 1ns/10ps

module and_tb;
    // Test signals
    reg clock_tb;
    reg clear_tb;
    reg PCout_tb, Zlowout_tb, MDRout_tb, R3out_tb, R7out_tb;
    reg MARin_tb, Zin_tb, PCin_tb, MDRin_tb, IRin_tb, Yin_tb;
    reg R3in_tb, R4in_tb, R7in_tb;
    reg [31:0] Mdatain_tb;
    wire [31:0] BusMuxOut_tb;

    // States for finite state machine
    parameter Default = 4'b0000, Reg_load1a = 4'b0001, Reg_load1b = 4'b0010, 
              Reg_load2a = 4'b0011, Reg_load2b = 4'b0100, 
              T0 = 4'b0101, T1 = 4'b0110, T2 = 4'b0111, T3 = 4'b1000, T4 = 4'b1001, T5 = 4'b1010;

    reg [3:0] Present_state = Default;

    // Instantiate the DataPath module
    DataPath DUT (
        .clock(clock_tb),
        .clear(clear_tb),
        .PCout(PCout_tb), .Zlowout(Zlowout_tb), .MDRout(MDRout_tb), 
        .R3out(R3out_tb), .R7out(R7out_tb),
        .MARin(MARin_tb), .Zin(Zin_tb), .PCin(PCin_tb), 
        .MDRin(MDRin_tb), .IRin(IRin_tb), .Yin(Yin_tb), 
        .R3in(R3in_tb), .R4in(R4in_tb), .R7in(R7in_tb),
        .Mdatain(Mdatain_tb),
        .BusMuxOut(BusMuxOut_tb),

        // Unconnected signals
        .R0out(), .R1out(), .R2out(), .R4out(), .R5out(), .R6out(), 
        .R8out(), .R9out(), .R10out(), .R11out(), .R12out(), .R13out(), 
        .R14out(), .R15out(), 
        .R0in(), .R1in(), .R2in(), .R5in(), .R6in(), .R8in(), .R9in(), 
        .R10in(), .R11in(), .R12in(), .R13in(), .R14in(), .R15in(),
        .HIin(), .HIout(), .LOin(), .LOout(), .Zhighout()
    );

    // Clock generation
    initial begin
        clock_tb = 0;
        forever #10 clock_tb = ~clock_tb;  // 10ns clock period
    end

    // FSM to control the states
    always @(posedge clock_tb) begin
        case (Present_state)
            Default: Present_state <= Reg_load1a;
            Reg_load1a: Present_state <= Reg_load1b;
            Reg_load1b: Present_state <= Reg_load2a;
            Reg_load2a: Present_state <= Reg_load2b;
            Reg_load2b: Present_state <= T0;
            T0: Present_state <= T1;
            T1: Present_state <= T2;
            T2: Present_state <= T3;
            T3: Present_state <= T4;
            T4: Present_state <= T5;
        endcase
    end

    // Control signal assignment based on the FSM states
    always @(Present_state) begin
        // Reset all signals to 0 by default
        PCout_tb = 0; Zlowout_tb = 0; MDRout_tb = 0;
        R3out_tb = 0; R7out_tb = 0; MARin_tb = 0; Zin_tb = 0;
        PCin_tb = 0; MDRin_tb = 0; IRin_tb = 0; Yin_tb = 0;
        R3in_tb = 0; R4in_tb = 0; R7in_tb = 0;
        Mdatain_tb = 32'h00000000;

        case (Present_state)
            Reg_load1a: begin  // Load value into R3
                Mdatain_tb <= 32'h00000022;
                MDRin_tb <= 1;
            end
            Reg_load1b: begin
                MDRin_tb <= 0;
                MDRout_tb <= 1; R3in_tb <= 1;
            end
            Reg_load2a: begin  // Load value into R7
                MDRout_tb <= 0; R3in_tb <= 0;
                Mdatain_tb <= 32'h00000024;
                MDRin_tb <= 1;
            end
            Reg_load2b: begin
                MDRin_tb <= 0;
                MDRout_tb <= 1; R7in_tb <= 1;
            end
            T0: begin
                MDRout_tb <= 0; R7in_tb <= 0;
                PCout_tb <= 1; MARin_tb <= 1;
            end
            T1: begin
                PCout_tb <= 0; MARin_tb <= 0;
                Mdatain_tb <= 32'h2A2B8000;  // Opcode for AND R4, R3, R7
                MDRin_tb <= 1;
            end
            T2: begin
                MDRin_tb <= 0;
                MDRout_tb <= 1; IRin_tb <= 1;
            end
            T3: begin
                MDRout_tb <= 0; IRin_tb <= 0;
                R3out_tb <= 1; Yin_tb <= 1;
            end
            T4: begin
                R3out_tb <= 0; Yin_tb <= 0;
                R7out_tb <= 1; Zin_tb <= 1;
            end
            T5: begin
                R7out_tb <= 0; Zin_tb <= 0;
                Zlowout_tb <= 1; R4in_tb <= 1;
            end
        endcase
    end

    // End simulation after some time
//    initial begin
//        #200 $finish;
//    end
endmodule
