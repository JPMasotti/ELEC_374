module outport(
input wire clk, clear, enable,
input wire [31:0] d,
output wire [31:0] q,

);